module LCD_1602(
				input              	CLK,               			// 50MHzʱ��
				input				RST_n,
				// Input frequency
				input	[71:0]		CLK_Data,	
				//LCD1602 Interface
				output             	LCD_EN,		// ʹ���ź�
				output 	reg         LCD_RS,     // ָ�����ѡ��
				output             	LCD_RW ,    // ����дѡ��
				output	reg	[7:0]	LCD_Data    // ��������
				);  

reg		[15:0] 		cnt;                         //������Ƶ�õ�lcd_clk
wire 				lcd_clk=cnt[15];     
reg 	[127:0] 	Line_Rom1 = "Frequency Count ";	//��ôд��wire��reg������
wire	[127:0]		Line_Rom2 = {"Data:",CLK_Data,"Hz"};


assign 	LCD_EN  = lcd_clk;                // ������ʱ�Ӹߵ�ƽ������                 
assign 	LCD_RW 	= 1'b0;                   // ֻд  

always @ (posedge CLK or negedge RST_n)
begin
	if(!RST_n)
		cnt <= 0;
	else
		cnt <= cnt + 1'b1;	
end
                                 
// ��������룺��40��״̬
parameter 	IDLE        	= 8'h00;	//���У���ʼ��
// дָ���ʼ��
parameter	DISP_SET     	= 8'h01;         // ��ʾģʽ����
parameter 	DISP_OFF     	= 8'h03;         // ��ʾ�ر�
parameter 	CLR_SCR      	= 8'h02;         // ��ʾ����
parameter 	CURSOR_SET1  	= 8'h06;         // ��ʾ����ƶ�����
parameter 	CURSOR_SET2  	= 8'h07;         // ��ʾ�����������
// ��ʾ��һ��
parameter 	ROW1_ADDR    	= 8'h05;         // д��1����ʼ��ַ
parameter 	ROW1_0       	= 8'h04;
parameter 	ROW1_1       	= 8'h0C;
parameter 	ROW1_2       	= 8'h0D;
parameter 	ROW1_3       	= 8'h0F;
parameter 	ROW1_4       	= 8'h0E;
parameter 	ROW1_5       	= 8'h0A;
parameter 	ROW1_6       	= 8'h0B;
parameter 	ROW1_7       	= 8'h09;
parameter 	ROW1_8       	= 8'h08;
parameter 	ROW1_9       	= 8'h18;
parameter 	ROW1_A       	= 8'h19;
parameter 	ROW1_B       	= 8'h1B;
parameter 	ROW1_C       	= 8'h1A;
parameter 	ROW1_D       	= 8'h1E;
parameter 	ROW1_E       	= 8'h1F;
parameter 	ROW1_F       	= 8'h1D;
// ��ʾ�ڶ���
parameter 	ROW2_ADDR    	= 8'h1C;         // д��2����ʼ��ַ
parameter 	ROW2_0       	= 8'h14;
parameter 	ROW2_1       	= 8'h15;
parameter 	ROW2_2       	= 8'h17;
parameter 	ROW2_3       	= 8'h16;
parameter 	ROW2_4       	= 8'h12;
parameter 	ROW2_5       	= 8'h13;
parameter 	ROW2_6       	= 8'h11;
parameter 	ROW2_7       	= 8'h10;
parameter 	ROW2_8       	= 8'h30;
parameter 	ROW2_9       	= 8'h31;
parameter 	ROW2_A       	= 8'h33;
parameter 	ROW2_B       	= 8'h32;
parameter 	ROW2_C       	= 8'h36;
parameter 	ROW2_D       	= 8'h37;
parameter 	ROW2_E       	= 8'h35;
parameter 	ROW2_F       	= 8'h34;

reg [5:0] current_state, next_state;    // ��̬����̬

// FSM: always1
always @ (posedge lcd_clk or negedge RST_n)
begin
	if(!RST_n)
		current_state <= IDLE;
	else
		current_state <= next_state;
end

// FSM: always2
always
begin
	case(current_state)
	IDLE        	: 	next_state = DISP_SET;
	// дָ���ʼ��
	DISP_SET    	: 	next_state = DISP_OFF;
	DISP_OFF    	: 	next_state = CLR_SCR;
	CLR_SCR     	:	next_state = CURSOR_SET1;
	CURSOR_SET1 	: 	next_state = CURSOR_SET2;
	CURSOR_SET2 	: 	next_state = ROW1_ADDR;
	// ��ʾ��һ��
	ROW1_ADDR   	: 	next_state = ROW1_0;
	ROW1_0      	: 	next_state = ROW1_1;
	ROW1_1      	: 	next_state = ROW1_2;
	ROW1_2      	: 	next_state = ROW1_3;
	ROW1_3      	: 	next_state = ROW1_4;
	ROW1_4      	: 	next_state = ROW1_5;
	ROW1_5      	: 	next_state = ROW1_6;
	ROW1_6      	: 	next_state = ROW1_7;
	ROW1_7      	: 	next_state = ROW1_8;
	ROW1_8      	: 	next_state = ROW1_9;
	ROW1_9      	: 	next_state = ROW1_A;
	ROW1_A      	: 	next_state = ROW1_B;
	ROW1_B      	: 	next_state = ROW1_C;
	ROW1_C      	: 	next_state = ROW1_D;
	ROW1_D      	: 	next_state = ROW1_E;
	ROW1_E      	: 	next_state = ROW1_F;
	ROW1_F      	: 	next_state = ROW2_ADDR;
	// ��ʾ�ڶ���
	ROW2_ADDR   	: 	next_state = ROW2_0; 
	ROW2_0      	: 	next_state = ROW2_1;
	ROW2_1      	: 	next_state = ROW2_2;
	ROW2_2      	: 	next_state = ROW2_3;
	ROW2_3      	:	next_state = ROW2_4;
	ROW2_4      	: 	next_state = ROW2_5;
	ROW2_5      	: 	next_state = ROW2_6;
	ROW2_6      	: 	next_state = ROW2_7;
	ROW2_7      	: 	next_state = ROW2_8;
	ROW2_8      	: 	next_state = ROW2_9;
	ROW2_9      	: 	next_state = ROW2_A;
	ROW2_A      	: 	next_state = ROW2_B;
	ROW2_B      	: 	next_state = ROW2_C;
	ROW2_C      	: 	next_state = ROW2_D;
	ROW2_D      	: 	next_state = ROW2_E;
	ROW2_E      	: 	next_state = ROW2_F;
	ROW2_F      	: 	next_state = ROW1_ADDR;
	default     	: 	next_state = IDLE ;
	endcase
end

// FSM: always3
always @ (posedge lcd_clk or negedge RST_n)
begin
	if(!RST_n)
		begin
		LCD_RS <= 0;
		LCD_Data <= 8'hxx;
		end
	else
		begin
			// дLCD_RS
			case(next_state)      
			IDLE        	: LCD_RS <= 0;	//ָ��
			// дָ���ʼ��
			DISP_SET    	: LCD_RS <= 0;	//ָ��
			DISP_OFF    	: LCD_RS <= 0;	//ָ��
			CLR_SCR     	: LCD_RS <= 0;	//ָ��
			CURSOR_SET1 	: LCD_RS <= 0;	//ָ��
			CURSOR_SET2 	: LCD_RS <= 0;	//ָ��
			// д���ݣ���ʾ��һ��
			ROW1_ADDR   	: LCD_RS <= 0;	//ָ��
			ROW1_0      	: LCD_RS <= 1;	//����
			ROW1_1      	: LCD_RS <= 1;	//����
			ROW1_2      	: LCD_RS <= 1;	//����
			ROW1_3      	: LCD_RS <= 1;	//����
			ROW1_4      	: LCD_RS <= 1;	//����
			ROW1_5      	: LCD_RS <= 1;	//����
			ROW1_6      	: LCD_RS <= 1;	//����
			ROW1_7      	: LCD_RS <= 1;	//����
			ROW1_8      	: LCD_RS <= 1;	//����
			ROW1_9      	: LCD_RS <= 1;	//����
			ROW1_A      	: LCD_RS <= 1;	//����
			ROW1_B      	: LCD_RS <= 1;	//����
			ROW1_C      	: LCD_RS <= 1;	//����
			ROW1_D      	: LCD_RS <= 1; 	//����
			ROW1_E      	: LCD_RS <= 1;	//����
			ROW1_F      	: LCD_RS <= 1;	//����
			// д���ݣ���ʾ�ڶ���
			ROW2_ADDR   	: LCD_RS <= 0;	//ָ��
			ROW2_0      	: LCD_RS <= 1;	//����
			ROW2_1     	: LCD_RS <= 1;	//����
			ROW2_2      	: LCD_RS <= 1;	//����
			ROW2_3      	: LCD_RS <= 1;	//����
			ROW2_4      	: LCD_RS <= 1;	//����
			ROW2_5      	: LCD_RS <= 1;	//����
			ROW2_6      	: LCD_RS <= 1;	//����
			ROW2_7      	: LCD_RS <= 1;	//����
			ROW2_8      	: LCD_RS <= 1;	//����
			ROW2_9      	: LCD_RS <= 1;	//����
			ROW2_A      	: LCD_RS <= 1;	//����
			ROW2_B      	: LCD_RS <= 1;	//����
			ROW2_C      	: LCD_RS <= 1;	//����
			ROW2_D      	: LCD_RS <= 1; 	//����
			ROW2_E      	: LCD_RS <= 1;	//����
			ROW2_F      	: LCD_RS <= 1;	//����
			endcase   

			// дLCD_Data
			case(next_state)
			IDLE        	: LCD_Data <= 8'hxx;
			// дָ���ʼ��
			DISP_SET    	: LCD_Data <= 8'h38;	//����16X2��ʾ,5X7����,8λ���ݽӿ�
			DISP_OFF    	: LCD_Data <= 8'h08;	//������ʾ���ܹ�,�޹��,����ʾ
			CLR_SCR     	: LCD_Data <= 8'h01;	//����ʾ,��긴λ��00Hλ��
			CURSOR_SET1 	: LCD_Data <= 8'h06;	//��ʾ��ַ��������дһ�����ݺ���ʾλ������һλ
			CURSOR_SET2 	: LCD_Data <= 8'h0C;	//������ʾ�����ع�꣬��겻��˸
			// д���ݣ���ʾ��һ��
			ROW1_ADDR   	: LCD_Data <= 8'h80;	//���ַ��ڵ�һ����ʾ
			ROW1_0      	: LCD_Data <= Line_Rom1[127:120];
			ROW1_1      	: LCD_Data <= Line_Rom1[119:112];
			ROW1_2      	: LCD_Data <= Line_Rom1[111:104];
			ROW1_3      	: LCD_Data <= Line_Rom1[103: 96];
			ROW1_4      	: LCD_Data <= Line_Rom1[ 95: 88];
			ROW1_5      	: LCD_Data <= Line_Rom1[ 87: 80];
			ROW1_6      	: LCD_Data <= Line_Rom1[ 79: 72];
			ROW1_7      	: LCD_Data <= Line_Rom1[ 71: 64];
			ROW1_8      	: LCD_Data <= Line_Rom1[ 63: 56];
			ROW1_9      	: LCD_Data <= Line_Rom1[ 55: 48];
			ROW1_A      	: LCD_Data <= Line_Rom1[ 47: 40];
			ROW1_B      	: LCD_Data <= Line_Rom1[ 39: 32];
			ROW1_C      	: LCD_Data <= Line_Rom1[ 31: 24];
			ROW1_D      	: LCD_Data <= Line_Rom1[ 23: 16]; 
			ROW1_E      	: LCD_Data <= Line_Rom1[ 15:  8];
			ROW1_F      	: LCD_Data <= Line_Rom1[  7:  0];
			// д���ݣ���ʾ�ڶ���
			ROW2_ADDR   	: LCD_Data <= 8'hC0;	//���ַ��ڵ�һ����ʾ
			ROW2_0      	: LCD_Data <= Line_Rom2[127:120];
			ROW2_1      	: LCD_Data <= Line_Rom2[119:112];
			ROW2_2      	: LCD_Data <= Line_Rom2[111:104];
			ROW2_3      	: LCD_Data <= Line_Rom2[103: 96];
			ROW2_4      	: LCD_Data <= Line_Rom2[ 95: 88];
			ROW2_5      	: LCD_Data <= Line_Rom2[ 87: 80];
			ROW2_6      	: LCD_Data <= Line_Rom2[ 79: 72];
			ROW2_7      	: LCD_Data <= Line_Rom2[ 71: 64];
			ROW2_8      	: LCD_Data <= Line_Rom2[ 63: 56];
			ROW2_9      	: LCD_Data <= Line_Rom2[ 55: 48];
			ROW2_A      	: LCD_Data <= Line_Rom2[ 47: 40];
			ROW2_B      	: LCD_Data <= Line_Rom2[ 39: 32];
			ROW2_C      	: LCD_Data <= Line_Rom2[ 31: 24];
			ROW2_D      	: LCD_Data <= Line_Rom2[ 23: 16];
			ROW2_E      	: LCD_Data <= Line_Rom2[ 15:  8];
			ROW2_F      	: LCD_Data <= Line_Rom2[  7:  0];
			endcase 
		end 
end

endmodule
